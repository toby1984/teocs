module not16(
input [15:0] in,
output [15:0] out);  

  not2 mynot0(in[ 0],out[0]); 
  not2 mynot1(in[ 1],out[1]); 
  not2 mynot2(in[ 2],out[2]); 
  not2 mynot3(in[ 3],out[3]); 
  not2 mynot4(in[ 4],out[4]); 
  not2 mynot5(in[ 5],out[5]); 
  not2 mynot6(in[ 6],out[6]); 
  not2 mynot7(in[ 7],out[7]); 
  not2 mynot8(in[ 8],out[8]); 
  not2 mynot9(in[ 9],out[9]); 
  not2 mynot10(in[10],out[10]); 
  not2 mynot11(in[11],out[11]);   
  not2 mynot12(in[12],out[12]);   
  not2 mynot13(in[13],out[13]);     
  not2 mynot14(in[14],out[14]);   
  not2 mynot15(in[15],out[15]);     
endmodule

module not2(input in,output out);  
  nand2 mynand(in,in,out); 
endmodule
